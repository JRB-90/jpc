`include "6502/CPU_6502.v"
`include "6522/VIA_6522.v"

module J6502_System (
    
);

VIA_6522 via1(

);

CPU_6502 cpu(

);

endmodule